module reservation_station (

  );

endmodule : reservation_station
