module pipeline_id (
  input clk,
  input rst,

  input [31:0] inst
  );

  

endmodule // pipeline_id
