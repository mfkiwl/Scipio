`include "common_def.h"

module exwb (
  input clk,
  input rst
  );

endmodule : exwb
