module id_reg_file;

endmodule // id_reg_file
